* SIMULATION
* -----------
.include "./sources/includes/32nm_HP.pm"

